`timescale 1ns/1ns
`include "Rsa256Core.sv"
`include "test/test_core.sv"
