`timescale 1ns/1ns
`include "utils/PipelineCtrl.v"
`include "utils/PipelineTb.v"
`include "Rsa256Core.sv"
`include "Rsa256Wrapper.sv"
`include "test/test_wrapper.sv"
